--  SALOME SALOMEDS : data structure of SALOME and sources of Salome data server 
--
--  Copyright (C) 2003  CEA/DEN, EDF R&D
--
--
--
--  File   : SALOMEDS_StudyPropertiesAttribute.cdl
--  Author : Yves FRICAUD
--  Module : SALOME

class StudyPropertiesAttribute from SALOMEDS inherits Attribute from TDF

	---Purpose: 


uses Attribute          from TDF,
     Label              from TDF,
     GUID               from Standard,
     DataSet            from TDF,
     RelocationTable    from TDF,
     Data               from TDF,
     ExtendedString     from TCollection,
     HSequenceOfExtendedString from TColStd,
     HSequenceOfInteger from TColStd

is    


    ---Purpose: class methods
    --          =============

    GetID (myclass)   
    ---C++: return const &  
    returns GUID from Standard;    

    Set (myclass; label : Label from TDF)
    returns StudyPropertiesAttribute from SALOMEDS;
    
    ---Purpose: Common methods
    --          ============
    
    Create 
    returns mutable StudyPropertiesAttribute from SALOMEDS;
    
    Init(me: mutable);

    SetUserName(me: mutable; theName : ExtendedString from TCollection);
    GetCreatorName(me) returns ExtendedString from TCollection;
    GetUserNames(me) returns HSequenceOfExtendedString from TColStd;
    SetFirstName(me: mutable; theName : ExtendedString from TCollection);
    
    SetModificationDate(me: mutable; theMinute, theHour, theDay, theMonth, theYear : Integer from Standard);
    GetCreationDate(me; theMinute, theHour, theDay, theMonth, theYear : out Integer from Standard)
    returns Boolean from Standard;
    GetModificationDates(me; theMinutes, theHours, theDays, theMonths, theYears : out HSequenceOfInteger from TColStd);
    
    SetCreationMode(me: mutable; theMode : Integer from Standard);
    GetCreationMode(me) returns Integer from Standard;

    SetModified(me: mutable; theModified : Integer from Standard);
    IsModified(me) returns Boolean from Standard;
    GetModified(me) returns Integer from Standard;
    
    SetLocked(me: mutable; theLocked : Boolean from Standard);
    IsLocked(me) returns Boolean from Standard;
    IsLockChanged(me: mutable; theErase : Boolean from Standard) returns Boolean from Standard;

    ID (me)
    	---C++: return const & 
    returns GUID from Standard;

    Restore (me: mutable; with : Attribute from TDF);

    NewEmpty (me)
    returns mutable Attribute from TDF;

    Paste (me; into : mutable Attribute from TDF;
	       RT   : mutable RelocationTable from TDF);

fields

    myUserName    : HSequenceOfExtendedString from TColStd;
    myMinute      : HSequenceOfInteger from TColStd;
    myHour        : HSequenceOfInteger from TColStd;
    myDay         : HSequenceOfInteger from TColStd;
    myMonth       : HSequenceOfInteger from TColStd;
    myYear        : HSequenceOfInteger from TColStd;
    myMode        : Integer from Standard;
    myModified    : Integer from Standard;
    myLocked      : Boolean from Standard;
    myLockChanged : Boolean from Standard;
    
end StudyPropertiesAttribute;
