//  File      : SALOMEDS_TargetAttribute.cdl
//  Created   : Fri Aug 16 10:20:05 2002
//  Author    : Yves FRICAUD
//  Project   : SALOME
//  Module    : SALOMEDS
//  Copyright : Open CASCADE 2002
//  $Header: 

class TargetAttribute from SALOMEDS inherits Relation from TDataStd

	---Purpose: 


uses Attribute         from TDF,
     Label             from TDF,
     GUID              from Standard,
     RelocationTable   from TDF,
     LabelList         from TDF

is    


    ---Purpose: class methods
    --          =============

    GetID (myclass)   
    ---C++: return const &  
    returns GUID from Standard;    

    Set (myclass; label : Label from TDF)
    returns TargetAttribute from SALOMEDS;
    
    ---Purpose: Comment methods
    --          ============
    
    Create 
    returns mutable TargetAttribute from SALOMEDS;
    
    Append(me: mutable; theReferencedObject : mutable Label form TDF);
    Get(me; theReferencedObjects : mutable : LabelList from TDF);
    Remove(me: mutable; theReferencedObject : mutable Label form TDF);

    ID (me)
    	---C++: return const & 
    returns GUID from Standard;

    Restore (me: mutable; with : Attribute from TDF);

    NewEmpty (me)
    returns mutable Attribute from TDF;

    Paste (me; into : mutable Attribute from TDF;
	       RT   : mutable RelocationTable from TDF);    

end TargetAttribute;
