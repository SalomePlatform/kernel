-- Copyright (C) 2005  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
-- CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
-- 
-- This library is free software; you can redistribute it and/or
-- modify it under the terms of the GNU Lesser General Public
-- License as published by the Free Software Foundation; either 
-- version 2.1 of the License.
-- 
-- This library is distributed in the hope that it will be useful 
-- but WITHOUT ANY WARRANTY; without even the implied warranty of 
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU 
-- Lesser General Public License for more details.
--
-- You should have received a copy of the GNU Lesser General Public  
-- License along with this library; if not, write to the Free Software 
-- Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
--
-- See http://www.salome-platform.org/ or email : webmaster.salome@opencascade.com
--
--
--
--  File   : SALOMEDS_PythonObjectAttribute.cdl
--  Author : Michael Ponikarov
--  Module : SALOME

class PythonObjectAttribute from SALOMEDS inherits Attribute from TDF

	---Purpose: 


uses Attribute          from TDF,
     Label              from TDF,
     GUID               from Standard,
     DataSet            from TDF,
     RelocationTable    from TDF,
     Data               from TDF,
     HArray1OfCharacter from TColStd

is    


    ---Purpose: class methods
    --          =============

    GetID (myclass)   
    ---C++: return const &  
    returns GUID from Standard;    

    Set (myclass; label : Label from TDF)
    returns PythonObjectAttribute from SALOMEDS;
    
    ---Purpose: Common methods
    --          ============
    
    Create 
    returns mutable PythonObjectAttribute from SALOMEDS;
    
    SetObject(me: mutable; theSequence : CString from Standard; theScript : Boolean from Standard);
    
    GetObject(me) returns CString from Standard;
    
    IsScript(me) returns Boolean from Standard;
    
    GetLength(me) returns Integer from Standard;

    ID (me)
    	---C++: return const & 
    returns GUID from Standard;

    Restore (me: mutable; with : Attribute from TDF);

    NewEmpty (me)
    returns mutable Attribute from TDF;

    Paste (me; into : mutable Attribute from TDF;
	       RT   : mutable RelocationTable from TDF);

fields

  mySequence : CString from Standard;
  myIsScript : Boolean from Standard;

end PythonObjectAttribute;
