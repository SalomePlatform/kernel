//  File      : SALOMEDS_SequenceOfRealAttribute.cdl
//  Created   : Wed Nov 28 16:20:40 2001
//  Author    : Yves FRICAUD
//  Project   : SALOME
//  Module    : SALOMEDS
//  Copyright : Open CASCADE 2001
//  $Header:



class SequenceOfRealAttribute from SALOMEDS inherits Attribute from TDF

	---Purpose: 


uses Attribute         from TDF,
     Label             from TDF,
     GUID              from Standard,
     HSequenceOfReal from TColStd,
     DataSet           from TDF,
     RelocationTable   from TDF,
     AttributeSequence from TDF,
     Data              from TDF,
     Comment           from TDataStd    	


is    


    ---Purpose: class methods
    --          =============

    GetID (myclass)   
    ---C++: return const &  
    returns GUID from Standard;    

    Set (myclass; label : Label from TDF)
    ---Purpose: Find, or create a Comment attribute and set the string.
    --          the Comment attribute is returned.
    returns SequenceOfRealAttribute from SALOMEDS;
    
    ---Purpose: Comment methods
    --          ============
    
    Create 
    returns mutable SequenceOfRealAttribute from SALOMEDS;
    
    ---Category: IntegerArray methods
    --          ===============

    Assign(me : mutable; other : HSequenceOfReal from TColStd);
    ---Purpose: Initialize the inner sequence by other one

    ChangeValue (me : mutable; Index : Integer from Standard; Value : Real);
    ---Purpose: Sets  the   <Index>th  element  of   the  sequence to <Value>
    
    Add (me : mutable; Value : Real from Standard);
    ---Purpose: Add  new value
    
    Value (me : mutable; Index : Integer from Standard) returns Real;
    ---Purpose: Value of index
    
    Remove (me : mutable; Index : Integer from Standard);
    ---Purpose: Remove element on index <Index>
 
    Length (me : mutable) returns Integer;
    ---Purpose: Returns length of sequence
 
    
    
    ID (me)
    	---C++: return const & 
    returns GUID from Standard;

    Restore (me: mutable; with : Attribute from TDF);

    NewEmpty (me)
    returns mutable Attribute from TDF;

    Paste (me; into : mutable Attribute from TDF;
	       RT   : mutable RelocationTable from TDF);    

fields

    myValue : HSequenceOfReal from TColStd;
    
end SequenceOfRealAttribute;
