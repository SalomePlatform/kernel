--  SALOME SALOMEDS : data structure of SALOME and sources of Salome data server 
--
--  Copyright (C) 2003  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
--  CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS 
-- 
--  This library is free software; you can redistribute it and/or 
--  modify it under the terms of the GNU Lesser General Public 
--  License as published by the Free Software Foundation; either 
--  version 2.1 of the License. 
-- 
--  This library is distributed in the hope that it will be useful, 
--  but WITHOUT ANY WARRANTY; without even the implied warranty of 
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU 
--  Lesser General Public License for more details. 
-- 
--  You should have received a copy of the GNU Lesser General Public 
--  License along with this library; if not, write to the Free Software 
--  Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA 
-- 
--  See http://www.opencascade.org/SALOME/ or email : webmaster.salome@opencascade.org 
--
--
--
--  File   : SALOMEDS_SequenceOfIntegerAttribute.cdl
--  Author : Yves FRICAUD
--  Module : SALOME

class SequenceOfIntegerAttribute from SALOMEDS inherits Attribute from TDF

	---Purpose: 


uses Attribute         from TDF,
     Label             from TDF,
     GUID              from Standard,
     HSequenceOfInteger from TColStd,
     DataSet           from TDF,
     RelocationTable   from TDF,
     AttributeSequence from TDF,
     Data              from TDF,
     Comment           from TDataStd    	


is    


    ---Purpose: class methods
    --          =============

    GetID (myclass)   
    ---C++: return const &  
    returns GUID from Standard;    

    Set (myclass; label : Label from TDF)
    ---Purpose: Find, or create a Comment attribute and set the string.
    --          the Comment attribute is returned.
    returns SequenceOfIntegerAttribute from SALOMEDS;
    
    ---Purpose: Comment methods
    --          ============
    
    Create 
    returns mutable SequenceOfIntegerAttribute from SALOMEDS;
    
    ---Category: IntegerArray methods
    --          ===============

    Assign(me : mutable; other : HSequenceOfInteger from TColStd);
    ---Purpose: Initialize the inner sequence by other one

    ChangeValue (me : mutable; Index, Value : Integer from Standard);
    ---Purpose: Sets  the   <Index>th  element  of   the  sequence to <Value>
    
    Add (me : mutable; value : Integer from Standard);
    ---Purpose: Add  new value
	
    Value (me : mutable; Index : Integer from Standard) returns Integer;
    ---Purpose: Value of index
     
    Remove (me : mutable; Index : Integer from Standard);
    ---Purpose: Remove element on index <Index>
 
    Length (me : mutable) returns Integer;
    ---Purpose: Returns length of sequence
 
    
    
    ID (me)
    	---C++: return const & 
    returns GUID from Standard;

    Restore (me: mutable; with : Attribute from TDF);

    NewEmpty (me)
    returns mutable Attribute from TDF;

    Paste (me; into : mutable Attribute from TDF;
	       RT   : mutable RelocationTable from TDF);    

fields

    myValue : HSequenceOfInteger from TColStd;
    
end SequenceOfIntegerAttribute;
