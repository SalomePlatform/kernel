-- Copyright (C) 2005  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
-- CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
-- 
-- This library is free software; you can redistribute it and/or
-- modify it under the terms of the GNU Lesser General Public
-- License as published by the Free Software Foundation; either 
-- version 2.1 of the License.
-- 
-- This library is distributed in the hope that it will be useful 
-- but WITHOUT ANY WARRANTY; without even the implied warranty of 
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU 
-- Lesser General Public License for more details.
--
-- You should have received a copy of the GNU Lesser General Public  
-- License along with this library; if not, write to the Free Software 
-- Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
--
-- See http://www.salome-platform.org/ or email : webmaster.salome@opencascade.com
--
--
--  File   : SALOMEDS_FileType.cdl
--  Author : Yves FRICAUD
--  Module : SALOME

class FileType from SALOMEDS inherits Comment from TDataStd

	---Purpose: 


uses Attribute         from TDF,
     Label             from TDF,
     GUID              from Standard,
     ExtendedString    from TCollection,
     DataSet           from TDF,
     RelocationTable   from TDF,
     AttributeSequence from TDF,
     Data              from TDF,
     Comment           from TDataStd


is    


    ---Purpose: class methods
    --          =============

    GetID (myclass)   
    ---C++: return const &  
    returns GUID from Standard;    

    Set (myclass; label : Label from TDF; 
	 Name : ExtendedString from TCollection)
    returns FileType from SALOMEDS;
    
    ---Purpose: Comment methods
    --          ============
    
    Create 
    returns mutable FileType from SALOMEDS;

    ID (me)
    	---C++: return const & 
    returns GUID from Standard;

    Restore (me: mutable; with : Attribute from TDF);

    NewEmpty (me)
    returns mutable Attribute from TDF;

    Paste (me; into : mutable Attribute from TDF;
	       RT   : mutable RelocationTable from TDF);    

end FileType;
