//  File      : SALOMEDS_TextHighlightColorAttribute.cdl
//  Created   : Wed Nov 28 16:20:40 2001
//  Author    : Yves FRICAUD
//  Project   : SALOME
//  Module    : SALOMEDS
//  Copyright : Open CASCADE 2001
//  $Header:




class TextHighlightColorAttribute from SALOMEDS inherits RealArray from TDataStd

	---Purpose: 


uses Attribute         from TDF,
     Label             from TDF,
     GUID              from Standard,
     ExtendedString    from TCollection,
     DataSet           from TDF,
     RelocationTable   from TDF,
     AttributeSequence from TDF,
     Data              from TDF,
     Comment           from TDataStd    	


is    


    ---Purpose: class methods
    --          =============

    GetID (myclass)   
    ---C++: return const &  
    returns GUID from Standard;    

    ---Purpose: Comment methods
    --          ============
    
    Create 
    returns mutable TextHighlightColorAttribute from SALOMEDS;

    ID (me)
    	---C++: return const & 
    returns GUID from Standard;

    Restore (me: mutable; with : Attribute from TDF);

    NewEmpty (me)
    returns mutable Attribute from TDF;

    Paste (me; into : mutable Attribute from TDF;
	       RT   : mutable RelocationTable from TDF);    

end TextHighlightColorAttribute;
